module And16_test;

    reg[15:0] a, b;
    wire[15:0] out;

    initial
        begin
            $dumpfile("And16_test.vcd");
            $dumpvars(0, and16);
            $monitor("a = %b, b = %b, out = %b", a, b, out);

            #1 a = 16'b0000000000000000; b = 16'b0000000000000000;
            #1 a = 16'b1111111111111111; b = 16'b1111111111111111;
            #1 a = 16'b0000000011111111; b = 16'b1111111100000000;
            #1 a = 16'b1111111100000000; b = 16'b0000000011111111;
            #1 a = 16'b0101010101010101; b = 16'b1010101010101010;
            #1 a = 16'b0000000011111111; b = 16'b0000000011111111;
            #1 a = 16'b1010101010101010; b = 16'b1010101010101010;
            #1 a = 16'b1111000011110000; b = 16'b1111000000001111;
            #1 $finish;
        end

    And16 and16(out, a, b);

endmodule

