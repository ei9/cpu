module Not16(out, in);

    output[15:0] out;
    input[15:0] in;

    Not not0(out[0], in[0]);
    Not not1(out[1], in[1]);
    Not not2(out[2], in[2]);
    Not not3(out[3], in[3]);
    Not not4(out[4], in[4]);
    Not not5(out[5], in[5]);
    Not not6(out[6], in[6]);
    Not not7(out[7], in[7]);
    Not not8(out[8], in[8]);
    Not not9(out[9], in[9]);
    Not not10(out[10], in[10]);
    Not not11(out[11], in[11]);
    Not not12(out[12], in[12]);
    Not not13(out[13], in[13]);
    Not not14(out[14], in[14]);
    Not not15(out[15], in[15]);

endmodule

